module top_module(
    output zero
);// Module body starts after semicolon
	assign zero = 0;
endmodule
